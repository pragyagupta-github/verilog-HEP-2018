module quiz(
reg[7:0]
