module adder(
input [15:0]a,b,
output [16:0]s);
assign s=a+b;
endmodule
