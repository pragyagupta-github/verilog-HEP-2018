module real_test;
real a;
initial
begin
a=12.22;
$display("a=%e",a);
end
endmodule
