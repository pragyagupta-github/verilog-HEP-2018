module grant(
input [3:0]a,
output out);

or a1(out,a[3],a[2],a[1],a[0]);
endmodule