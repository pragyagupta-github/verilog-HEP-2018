// 4*4  multiplier
module multiplier(
input [3:0]x,y,
output [7:0]out);
wire [21:0]w;
wire [10:0]c;

and g1(out[0], x[0], y[0]),
    g2(w[0], x[1], y[0]),
    g3(w[1], x[2], y[0]),
    g4(w[2], x[3], y[0]),

    g5(w[3], x[0], y[1]),
    g6(w[4], x[1], y[1]),
    g7(w[5], x[2], y[1]),
    g8(w[6], x[3], y[1]),

    g9(w[7], x[0], y[2]),
    g10(w[8], x[1], y[2]),
    g11(w[9], x[2], y[2]),
    g12(w[10], x[3], y[2]),

    g13(w[11], x[0], y[3]),
    g14(w[12], x[1], y[3]),
    g15(w[13], x[2], y[3]),
    g16(w[14], x[3], y[3]);

fulladder_ha f1(w[3],w[0],1'b0,out[1],c[0]),
             f2(w[4],w[1],c[0],w[8],c[1]),
             f3(w[5],w[2],c[1],w[9],c[2]),
             f4(w[6],1'b0,c[2],w[10],c[3]),

             f5(w[11],w[8],1'b0,out[2],c[4]),
             f6(w[12],w[9],c[4],w[15],c[5]),
             f7(w[13],w[10],c[5],w[16],c[6]),
             f8(w[14],c[3],c[6],w[17],c[7]),

             f9(w[18],w[15],1'b0,out[3],c[8]),
             f10(w[19],w[16],c[8],out[4],c[9]),
             f11(w[20],w[17],c[9],out[5],c[10]),
             f12(w[21],c[10],c[7],out[6],out[7]);

endmodule
